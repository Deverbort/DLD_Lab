library verilog;
use verilog.vl_types.all;
entity OP_TB is
end OP_TB;
